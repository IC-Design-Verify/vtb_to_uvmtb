// ***********************************************************************
// *****************                                                       
// ***** ***********                                                       
// *****   *********                                                       
// *****     *******      Copyright (c) 2025  Kang Yaopeng  
// *****       *****                                                       
// *****     *******             All rights reserved                       
// *****   *********                                                       
// ***** ***********                                                       
// *****************                                                       
// ***********************************************************************
// PROJECT        : 
// FILENAME       : ahb_agent_pkg.sv
// Author         : IC_VERIFY
// LAST MODIFIED  : 2025-09-10 13:53
// ***********************************************************************
// DESCRIPTION    :
// ***********************************************************************
// $Revision: $
// $Id: $
// ***********************************************************************
package ahb_agent_pkg;
  import uvm_pkg::*;

  `include "ahb_driver.svh"
endpackage
// ***********************************************************************
// $Log: $
// $Revision $

// ***********************************************************************
// *****************                                                       
// ***** ***********                                                       
// *****   *********                                                       
// *****     *******      Copyright (c) 2025  Kang Yaopeng  
// *****       *****                                                       
// *****     *******             All rights reserved                       
// *****   *********                                                       
// ***** ***********                                                       
// *****************                                                       
// ***********************************************************************
// PROJECT        : 
// FILENAME       : ahb_intf.sv
// Author         : yaopeng.kang
// LAST MODIFIED  : 2025-09-06 16:37
// ***********************************************************************
// DESCRIPTION    :
// ***********************************************************************
// $Revision: $
// $Id: $
// ***********************************************************************
interface ahb_intf(input bit hclk, 
                   input bit hrst_n);

  logic[31:0] haddr ;
  logic[3 :0] hprot ;
  logic[31:0] hrdata;
  logic[0 :0] hready;
  logic[1 :0] hresp ;
  logic[0 :0] hsel  ;
  logic[1 :0] htrans;
  logic[31:0] hwdata;
  logic[0 :0] hwrite;


endinterface
// ***********************************************************************
// $Log: $
// $Revision $
